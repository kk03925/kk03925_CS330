module Adder
(
	input [63:0] a,
	input [63:0] b,
	
	output reg [63:0] out
);

	always@(a or b)
		begin
			out = a+b;
		end
endmodule