module tb
(




);

	
	initial
	clk = 1'b0;
	
	always
	#5 clk = ~clk;
	
	initial
	begin
		
	
	
	
	end